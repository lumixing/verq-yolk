module verq

pub struct User {
pub:
	username string
	id       string
}
